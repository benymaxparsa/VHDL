-- A General Purpose Shift Register with Shift-to-left, Shift-to-right, Reset, and Counter abilities 

